module hello;
    initial
    begin
        $display("Hello bich!");
        $finish;
    end
endmodule