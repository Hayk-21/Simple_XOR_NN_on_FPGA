module my_xor(input logic signed [31:0] x, output reg signed [31:0] pred);

endmodule